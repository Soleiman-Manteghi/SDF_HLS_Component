// SDF_HLS_componentqsys_component_0.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module SDF_HLS_componentqsys_component_0 (
		input  wire        clock,    // clock.clk
		input  wire        resetn,   // reset.reset_n
		input  wire [31:0] s0_data,  //    s0.data
		output wire        s0_ready, //      .ready
		input  wire        s0_valid, //      .valid
		output wire [31:0] s4_data,  //    s4.data
		input  wire        s4_ready, //      .ready
		output wire        s4_valid  //      .valid
	);

	SDF_HLS_component_internal sdf_hls_component_internal_inst (
		.clock    (clock),    // clock.clk
		.resetn   (resetn),   // reset.reset_n
		.s0_data  (s0_data),  //    s0.data
		.s0_ready (s0_ready), //      .ready
		.s0_valid (s0_valid), //      .valid
		.s4_data  (s4_data),  //    s4.data
		.s4_ready (s4_ready), //      .ready
		.s4_valid (s4_valid)  //      .valid
	);

endmodule
